AC-PHASE-SHIFT
V1 1 0 SIN(0 1 60)
R1 1 2 1
R2 1 3 1
L1 2 0 1
R3 3 0 6.3E3
.TRAN 2.5E-3 4E-2 0
.PROBE
.END