EG16.35
V1 1 0 AC 1E-3
RCC 1 2 1E3
CC1 2 3 1E-6
RB1 6 3 90E3
RB2 3 0 10E3
RC 6 4 5E3
RE 5 0 1E3
CB 5 0 4.7E-6
CC2 4 7 4.7E-6
RL 7 0 5E3
VCC 6 0 DC 20
Q 4 3 5 Q2N2222
.LIB EVAL.LIB
.AC DEC 100 10 10E6
.PROBE
.END