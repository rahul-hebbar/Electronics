EG16.24
VCC 5 0 DC 5
V1 1 0
R1 5 2 5E3
R2 5 4 2E3
R3 5 7 100
R4 5 10 5E3
R5 6 0 1E3
Q1 3 2 1 Q2N3904
Q2 4 3 6 Q2N3904
Q4 7 4 8 Q2N3904
Q3 9 6 0 Q2N3904
Q5 11 10 9 Q2N3904
D1 8 9 D1N4148
D2 11 12 D1N4148
D3 12 0 D1N4148
.LIB EVAL.LIB
.DC V1 0 5 0.01
.TF V(9) V1
.PROBE
.END