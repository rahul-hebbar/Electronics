FULL-WAVE-BRIDGE-RECTIFER
V1 1 0 SIN(0 15 60)
D1 1 2 DMOD
D3 3 1 DMOD
D2 0 2 DMOD
D4 3 0 DMOD
RL 2 3 10E3
*CL 2 3 3.5E-6
.MODEL DMOD D 
.TRAN 2.5E-3 5E-2 0
.PROBE V(2,3)
.END