NON-INV-OPAMP
R2 1 0 10E3
R1 1 3 20E3
R3 2 0 10E3
V1 2 0 DC 5
E1 3 0 2 1 999E3
.DC V1 5 5 1
.PRINT DC V(3)
.END