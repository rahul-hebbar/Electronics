EG8.3
C1 1 0 0.1 IC=9
R1 1 0 9
S1 1 2 5 0 SMOD
S2 1 3 6 0 SMOD
R2 2 0 4.5
R3 3 0 72
.MODEL SMOD VSWITCH (VT=0.5)
V0 5 0 PWL(0 0 1 0 1 1)
V1 6 0 PWL(0 1 1 1 1 0)
.TRAN 0.01 2 UIC
.PROBE
.END
