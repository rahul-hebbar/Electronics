eg16.15
V1 1 0 AC 1
C1 1 2 0.16E-6
R1 2 0 1E3
.AC LIN 100 1 5000
.PROBE
.END