EG16.10
V1 1 0 PWL(0 0 0.001 1 15 1)
R 1 2 2
C 2 0 2
.TRAN 0.1 15 0
.PROBE
.END