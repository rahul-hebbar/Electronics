INST-OPAMP
V1 1 0 DC 0
RB1 1 0 10E3
V2 4 0 DC 5
RB2 4 0 10E3
R1 3 2 10E3
R2 5 6 10E3
RG 2 5 10E3
R3 3 7 10E3
R5 6 8 10E3
R6 8 0 10E3
R4 7 9 10E3
RL 9 0 10E3
E1 3 0 1 2 999E3
E2 6 0 4 5 999E3
E3 9 0 8 7 999E3
.DC V1 0 10 0.1
.PROBE
.END