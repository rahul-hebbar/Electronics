EG1 MULTIDCSOURCE
V1 1 0 DC 24
R1 1 2 10E3
R2 2 3 8.1E3
R3 2 0 4.7E3
V2 3 0 DC 15
.END