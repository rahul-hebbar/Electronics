EG16.28
VGS 1 0
VDS 2 0
M 2 1 0 0 IRF150
.LIB EVAL.LIB
.DC VDS 0 1 0.01 VGS 2.8 3.3 0.1
.PROBE
.END