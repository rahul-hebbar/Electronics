EG16.32
VCC 5 0 DC 10V
RC 5 2 980
RB1 5 3 26E3
RB2 3 0 26E3
RE 4 0 2E3
CC 1 3 10E-6
Q 2 3 4 QMOD
.MODEL QMOD NPN (IS=3.6E-15)
V1 1 0 AC 1E-6
.AC LIN 1000 1 1E4
.PROBE
.END