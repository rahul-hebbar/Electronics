eg16.6
V1 1 0 DC 0.1
R1 1 2 1E3
R2 2 4 20E3
R3 3 0 1E3
R4 3 4 10E3
E1 4 0 3 2 1G
.END