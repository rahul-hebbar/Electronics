EG16.21
V1 1 0 DC 10
R1 1 2 2.7E3
R2 1 3 330E3
R3 4 0 1E3
Q1 2 3 4 QMOD
.MODEL QMOD NPN (IS=3.9E-15)
.OP
.END