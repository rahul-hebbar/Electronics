INVERTER_RESISTIVE_LOAD
V1 1 0 DC 1
VDD 3 0 DC 10
R1 3 2 2E3
M1 2 1 0 0 NMOD
.MODEL NMOD NMOS (KP=0.5E-3 VTO=1)
.DC V1 0 10 0.01
.PROBE
.END