EG16.27
V1 1 0 DC 12
M1 1 1 2 2 NMOD
M2 2 3 0 0 NMOD
VG 3 0 DC 12
.MODEL NMOD NMOS (KP=0.5E-3 VTO=2)
.OP
.END