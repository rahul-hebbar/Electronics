eg16.4
V1 1 0 DC 3
R1 1 2 2
R2 2 0 6
R3 2 3 1
R4 3 0 8
G1 3 0 2 0 0.25
.OP
.END