EG16.23
IB 0 1
VCE 2 0
Q 2 1 0 Q2N3904
.LIB EVAL.LIB
.DC VCE 0 5 0.1 IB 0 20E-6 4E-6
.PROBE
.END