SEDRA5.10
VDD 1 0 DC 15
RD 1 2 10E3
M1 2 3 0 0 NMOD
RGD 2 3 10E6
CC1 5 3 1E-6
VIN 5 0 AC 1E-6
CC2 2 4 1E-6
RL 4 0 10E3
.MODEL NMOD NMOS (KP=0.25E-3 VTO=1.5 LAMBDA=0.02)
.AC DEC 1000 1 1E6
.OP
.PROBE
.END