ACSINE
V1 1 0 SIN(0 15 60)
R1 1 0 10E3
.TRAN 2E-3 20E-3 0
.PROBE
.END