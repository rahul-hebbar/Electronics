TEST2
VDD 3 0 DC 10
RD 3 2 1E3
M1 2 1 0 0 NMOD
.MODEL NMOD NMOS (KP=10E-3 VTO=2)
VG 1 0 4
C1 2 0 100E-12 IC=10
.TRAN 10E-9 400E-9
.PROBE
.END