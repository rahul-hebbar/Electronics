EG8.4
C1 1 0 0.25 IC=10
R1 1 0 4
G 0 1 1 0 0.75
.TRAN 0.01 2 UIC
.PROBE
.END