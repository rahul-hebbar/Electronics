EG16.22
VB 1 0 DC 5
RB 1 3 20E3
VCC 4 0 DC 5
RC 4 2 1E3
D 3 2 DMOD
.MODEL DMOD D (IS=2.3E-11)
Q 2 3 0 BMOD
.MODEL BMOD npn (IS=8.75E-15 BF=50)
.OP
.END