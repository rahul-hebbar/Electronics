eg16.5
V1 1 0 DC 1
V2 1 2 0
R1 2 3 150
R2 3 0 25
R4 4 0 1.5E3
R3 1 4 15E3
F1 4 3 V2 50
.op
.end