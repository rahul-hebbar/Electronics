LOW-PASS-FILTER
V2 1 0 DC 24
V1 2 1 AC 24
L1 2 3 100E-3
L2 3 4 250E-3
C1 3 0 100E-6
RL 4 0 1E3
.AC LIN 30 500 15E3
.PRINT AC V(4)
.PROBE
.END