eg16.13
V1 1 0 AC 6 -90
R1 1 2 1
C1 2 0 0.5
.AC LIN 1 0.31831 0.31831
.PRINT AC VM(C1) VP(C1) IM(C1) IP(C1)
.END