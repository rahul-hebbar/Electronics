EG16.25
V1 1 0 DC 18
RD 1 2 500
RS 3 0 1000
J 2 0 3 JMOD
.MODEL JMOD NJF (BETA=0.5E-3 VTO=-4)
.OP
.END