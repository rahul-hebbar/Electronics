TRANSIENT_1
V1 1 0 PWL(0 12 40 12 40 24)
R1 1 2 6E3
R2 3 0 3E3
C1 2 0 0.5E-3 IC=0
*SWITCH INPUT
V2 4 0 PWL(0 -1 50 -1 50 1)
R3 4 0 1
*MODEL VOLTAGE CONTROLLED SWITCH
S1 2 3 4 0 SMOD
.MODEL SMOD VSWITCH (VT=0)
.TRAN 0.01 100 0 UIC
.OP
.PROBE
.END