TEST1
VGS 1 0
VDS 2 0
M1 2 1 0 0 NMOD
.MODEL NMOD NMOS (KP=0.5E-3 VTO=2)
.DC VDS 0 2 0.01 VGS 1.8 3 0.2
.PROBE
.END