eg16.12
V1 1 0 EXP(0 10 1 10 50 10)
R1 1 0 1
.TRAN 0.01 100 0
.PROBE
.END