PD_FWBR_V_CHAR
*V1 1 0 DC 1
V1 1 0 SIN(0 4 1)
R1 1 2 1E3
R2 2 3 2E3
E1 4 0 0 2 1E9
R3 2 5 2E3
D1 3 4 DMOD
D2 4 5 DMOD
R4 3 6 2E3
R5 6 7 2E3
E2 7 0 5 6 1E9
.MODEL DMOD D
*.DC V1 -5 5 0.05
.TRAN 0.01 2 0
.PROBE V(7) V(1)
.END