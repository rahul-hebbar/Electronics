LOW-PASS-FILTER
V1 1 0 AC 10
R1 1 2 680
L1 2 3 108E-3
L2 3 4 108E-3
C1 3 0 0.47E-6
R2 4 0 680
.AC LIN 100 1 5000
.PROBE
.END