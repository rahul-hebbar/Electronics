OPAMP
V1 1 0 DC 0.1
R1 1 3 1E3
R2 2 0 1E3
R3 2 6 100E3
RL 6 0 10E3
XOPAMP 3 2 7 4 6 uA741
VS1 7 0 DC 15
VS2 4 0 DC -15
.LIB EVAL.LIB
.TRAN 1 1
.PRINT TRAN V(6)
.END