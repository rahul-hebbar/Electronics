CS_MULTISTAGE
VSIG 1 8 AC 1E-3
VBIAS 8 0 DC 2
RIN 1 2 200
VDD 5 0 12
RD1 5 4 1E3
M1 4 2 3 3 NMOD1
RS 3 0 200
CBY 3 0 500E-9
CB 4 6 100E-9
RVB1 5 6 100E3
RVB2 6 0 10E3
RD2 5 7 1E3
M2 7 6 0 0 NMOD2 
.MODEL NMOD1 NMOS (CGSO=250E-12 CGDO=80E-12 VTO=1 KP=0.02)
.MODEL NMOD2 NMOS (CGSO=250E-12 CGDO=80E-12 VTO=0.5 KP=0.115)
.OP
.PROBE
.AC DEC 1000 1 1E10
.END