TRANSIENT_2
V1 1 0 PULSE(1 0 10m 0.1u 0.1u 10m 20m)
R1 2 1 10E3
C1 2 0 1E-6 IC=0
.TRAN 1m 100m 0 UIC
.PROBE
.END