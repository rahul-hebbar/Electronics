EG16.30
VDD 3 0 DC 12
VGG 1 0
M1 2 1 0 0 NMOD
.MODEL NMOD NMOS (KP=0.5E-3 VTO=2)
M2 3 3 2 2 PMOD
.MODEL PMOD PMOS (KP=0.5E-3 VTO=-2)
.DC VGG 0 12 0.05 NMOS NMOD(KP) 0.5E-3 0.1E-3 0.4E-3
.PROBE
.END 