eg16.2
V1 1 0 DC 24
R1 1 2 2
R2 2 0 6
V2 2 3 DC 4
R3 3 0 8
I1 3 0 DC 3
.END