V_CHAR_CLIPPER
V1 1 0 DC 1
E 4 0 1 2 1E9
R1 2 4 10
D1 3 2 DMOD
D2 3 0 DMOD
.MODEL DMOD D(IS=10E-9 N=2 BV=5)
.DC V1 -15 15 0.1
.PROBE V(2)
.END