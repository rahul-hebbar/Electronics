EG16.16
V1 1 0 AC 1
R1 1 2 1E3
C1 2 0 0.16E-6
.AC DEC 100 1 100E3
.PROBE
.END