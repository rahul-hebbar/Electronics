EG16.26
V1 1 0 DC 12
M1 1 1 2 2 NMOD
M2 2 0 0 0 NMOD
.MODEL NMOD NMOS (VTO=-4 KP=2E-3)\
.OP
.END