OPAMP_SELF
V1 1 0 DC 0.1
R1 1 3 1E3
R2 2 0 1E3
R3 2 6 100E3
RL 6 0 10E3
E 6 0 3 2 10E6
.TRAN 1 1
.PRINT TRAN V(6)
.END