MOS_FB_AMP
VS 1 0 AC 1E-6
C1 1 2 10E-6
RF 2 3 1E6
RD 4 3 4E3
C2 3 5 10E-6
RL 5 0 6E3
VDD 4 0 DC 22
M1 3 2 0 0 NMOD
.MODEL NMOD NMOS (KP=0.5E-3 VTO=2)
.AC LIN 1 100E3 100E3
.PRINT AC VM(5) VM(1) VP(5)
.PROBE
.TF V(3) VS
.OP
.END