eg16.3
V1 1 0 DC 5
R1 1 2 2
R2 2 0 1
R3 2 4 5
R4 4 3 3
R5 4 0 4
E1 0 3 2 0 10
.OP
.END