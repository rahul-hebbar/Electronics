eg16.1
V1 3 0 DC 28
R1 3 1 5
R2 1 0 4
R3 1 2 1
R4 2 0 3
.END