eg16.34
V1 1 0 AC 1
R4 6 0 4E3
R1 1 2 1E3
R2 3 4 1E6
R3 5 4 1E3
C1 2 3 10E-6
C2 4 6 10E-6
V2 5 0 DC 10
M1 4 3 0 0 MMOD
.MODEL MMOD NMOS (VTO=2 KP=0.5E-3 CGSO=10E-6 )
.AC DEC 100 1 10E5
.PRINT AC VP(6) V(3)
.TF V(4) V1
.OP
.PROBE
.END
