EG16.20
V1 1 0 SIN(0 24 60)
D1 1 2 D1N4148
C1 2 0 10E-6
R1 2 0 10E3
.LIB EVAL.LIB
.TRAN 2E-6 50E-3 0
.PROBE
.END