INV-OPAMP
V1 2 0 DC 0
R1 2 1 1.18E3
R2 1 3 3.29E3
E1 3 0 0 1 999E3
.DC V1 3.5 0 0.1
.PROBE
.END