AC-RES-CAP
V1 1 0 SIN(0 0.5 60)
R1 1 2 30
C1 2 0 100E-6
.TRAN 0.025 0.05 0
.PROBE
.END