eg16.17
V1 1 0 DC 3
R1 2 0 1E3
D1 1 2 DMOD
.MODEL DMOD D (Is=10e-9 N=2)
.TEMP 300
.OP
.END