eg16.19
V1 1 0 SIN(0 24 1)
R1 1 2 1E3
D1 2 3 DMOD
D2 0 3 DMOD
.MODEL DMOD D (IS=10E-9 N=2 BV=12)
.TRAN 0.01 2
.PROBE
.END