EG8.5
V1 1 0 10
R1 1 2 5
L1 2 0 2 IC=1
.TRAN 0.01 3 UIC
.PROBE
.END