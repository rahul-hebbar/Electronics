MULTI-AC-SRC
V1 1 0 AC 55
V2 4 0 AC 43 25
L1 1 2 450E-3
L2 2 3 150E-3
R1 3 4 1E-12
C1 2 0 330E-6
.AC LIN 1 30 30
.PRINT AC V(2,0)
.END