DIODE_FWBR_V_CHAR
V1 1 0 DC 1
D1 1 2 DMOD
D3 3 1 DMOD
D2 0 2 DMOD
D4 3 0 DMOD
RL 2 3 10E3
.MODEL DMOD D
.DC V1 -10 10 0.1
.PROBE V(2,3)
.OP
.END