OPAMP-INT-SQ-INP
VIN 1 0 PULSE(0 1 0 1E-9 1E-9 0.001 0.002)
R1 2 1 100
C1 2 3 100E-8
R2 2 3 200
.SUBCKT OPAMP 1 2 3 4
E1 1 2 3 4 999E3
.ENDS
X1 3 0 0 2 OPAMP
.TRAN 0.001 0.01 0
.PROBE
.END