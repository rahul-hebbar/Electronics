EG16.36
R1 1 5 6.5E3
R2 1 2 188.5E3
C1 3 2 1E-9 IC=5
C2 4 3 1E-9
C3 5 4 1E-9
R3 3 0 6.5E3
R4 4 0 6.5E3
E 2 0 0 1 10E6
.TRAN 1E-6 800E-6 UIC
.PROBE
.END 