OPAMP-INT-SIN-INP
VIN 1 0 SIN(0 1 50)
R1 2 1 100
C1 2 3 100E-8
R2 2 3 200
E1 3 0 0 2 999E3
.TRAN 0.01 50E-3 0
.PROBE
.END