EG2.2
V1 1 0 SIN(0 6 0.159 0 0 90)
R1 1 0 1
R2 1 0 2
R3 1 0 3
.TRAN 0.1 10
.PROBE
.END
