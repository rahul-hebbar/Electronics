EG16.29
VDD 3 0 DC 12
M1 2 1 3 3 PMOD
M2 2 1 0 0 NMOD
.MODEL PMOD PMOS (KP=0.5E-3 VTO=-2)
.MODEL NMOD NMOS (KP=0.5E-3 VTO=2)
VG 1 0
.DC VG 0 12 0.01
.PROBE
.END
