EG8.2
R1 1 0 5
S1 1 2 6 0 SMOD
R2 2 0 20
L1 2 0 8 IC=10
VC 6 0 PWL(0 0 0.4 0 0.4 1)
.MODEL SMOD VSWITCH (VT=0.5)
.TRAN 0.01 1.4
.PROBE
.END