eg16.9
R1 1 0 2
L1 1 2 1 IC=-0.32
C1 2 0 0.02 IC=2
.TRAN 0.05 3 0 UIC
.PROBE
.END