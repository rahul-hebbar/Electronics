TEST3_CSAMP_SELF
V1 1 0 AC 1E-3
CC1 1 2 1E-6
RB1 3 2 2E6
RB2 2 0 1E6
VD 3 0 12
RD 3 4 4E3
CC2 4 5 1E-6
RL 5 0 4E3
M1 4 2 0 0 NMOD
.MODEL NMOD NMOS (KP=0.5E-3 VTO=2)
.AC DEC 1000 1 1E6
.PROBE
.END