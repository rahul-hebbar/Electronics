RCCKT
V1 1 0 DC 10
C1 1 2 47E-6 IC=0
C2 1 2 22E-6 IC=0
R1 2 0 3.3E3
.TRAN 0.01 2 0
.PROBE
.END