EG16.11
V1 1 0 PULSE(0 1 0 0.001)
R1 1 2 1
L1 2 0 4
C1 2 0 1
.TRAN 0.01 10 0
.PROBE
.END